module Shifter( result, leftRight, shamt, sftSrc  );
    
  output wire[31:0] result;

  input wire leftRight;
  input wire[4:0] shamt;
  input wire[31:0] sftSrc ;
  
  assign result=(leftRight==1)? sftSrc<<shamt:sftSrc>>shamt;
  /*your code here*/ 
	
endmodule